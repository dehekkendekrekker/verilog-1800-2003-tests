//----------------------------------------------------------------
// Tests support of simple_immediate_assertions: assert()
//----------------------------------------------------------------
module simple_immediate_assert_statement();

initial assert(0);

endmodule
